library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity ch4_ROM is
    Port (
        ROMaddress : in integer range 0 to 65535;        -- ROM access address
        
        sub_ch1_vec : out std_logic_vector(20 downto 0); -- sub channel-1 input vector
        sub_ch2_vec : out std_logic_vector(20 downto 0); -- sub channel-2 input vector
        sub_ch3_vec : out std_logic_vector(20 downto 0); -- sub channel-3 input vector
        sub_ch4_vec : out std_logic_vector(20 downto 0)  -- sub channel-4 input vector
    );
end ch4_ROM;

architecture Behavioral of ch4_ROM is
    type ROM_entry is array (0 to 3) of std_logic_vector(20 downto 0);
    type ROM_type is array (0 to 289) of ROM_entry;
    signal ch_ROM : ROM_type := ( 
    ("000000000000000000000",	"000000000000000000000",	"000000000000000000000",	"000000000000000000000"),
    ("110000001000011111111",	"000000000000000000000",	"000000000000000000000",	"000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001111101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001111101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001111101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001011001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001100011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001101001111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000111111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001010011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000010000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001000011111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("110000001110101111111",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000"),
    ("000000000000000000000",    "000000000000000000000",    "000000000000000000000",    "000000000000000000000")
    );

begin

    sub_ch1_vec <= ch_ROM(ROMaddress)(0);
    sub_ch2_vec <= ch_ROM(ROMaddress)(1);
    sub_ch3_vec <= ch_ROM(ROMaddress)(2);
    sub_ch4_vec <= ch_ROM(ROMaddress)(3);

end Behavioral;