library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity ch2_timer_ROM is
    Port (
        reset_time : in std_logic;                      -- reset time counter to 0 
        tempo_clock: in std_logic;                      -- 100MHz clock for timer signal update counter
        
        ROMaddress : out integer range 0 to 65535;      -- global timing signal
        checker_s  : out std_logic
    );
end ch2_timer_ROM;

architecture Behavioral of ch2_timer_ROM is
    type ROM_type is array (0 to 170) of std_logic_vector(20 downto 0);
    signal time_ROM : ROM_type := (
    "000000000000000000000",
    "000000000000000000000",
    "000001101010111000000",
    "000001101100110000000",
    "000001101110101000000",
    "000001110000000010000",
    "000001110011110010000",
    "000001110110100110000",
    "000001110111000100000",
    "000001110111100010000",
    "000001111000011110000",
    "000001111000111100000",
    "000001111001011010000",
    "000001111001111000000",
    "000001111010010110000",
    "000001111010110100000",
    "000001111011010010000",
    "000001111011110000000",
    "000001111100001110000",
    "000001111100101100000",
    "000001111101001010000",
    "000001111101101000000",
    "000001111110000110000",
    "000001111110100100000",
    "000001111111000010000",
    "000010000010110010000",
    "000010000100101010000",
    "000010000110100010000",
    "000010001000111000000",
    "000010001010110000000",
    "000010001100101000000",
    "000010001110000010000",
    "000010010000011000000",
    "000010010001110010000",
    "000010010100001000000",
    "000010010100100110000",
    "000010010101000100000",
    "000010010101100010000",
    "000010010110011110000",
    "000010010110111100000",
    "000010010111011010000",
    "000010010111111000000",
    "000010011000010110000",
    "000010011000110100000",
    "000010011001010010000",
    "000010011001110000000",
    "000010011010001110000",
    "000010011010101100000",
    "000010011011001010000",
    "000010011011101000000",
    "000010011100000110000",
    "000010011100100100000",
    "000010011101000010000",
    "000010011101100000000",
    "000010011101110100000",
    "000010011110001000000",
    "000010011110011100000",
    "000010011110110000000",
    "000010011111000100000",
    "000010011111011000000",
    "000010011111101100000",
    "000010100000000000000",
    "000010100000010100000",
    "000010100000101000000",
    "000010100000111100000",
    "000010100001010000000",
    "000010100100100010000",
    "000010100101000000000",
    "000010100101111100000",
    "000010101010101000000",
    "000010101100000010000",
    "000010110000010000000",
    "000010110010001000000",
    "000010110011100010000",
    "000010110101111000000",
    "000010110110010110000",
    "000010110110110100000",
    "000010110111010010000",
    "000010110111110000000",
    "000010111011000010000",
    "000010111101011000000",
    "000010111110110010000",
    "000011000010000100000",
    "000011000010011000000",
    "000011000010101100000",
    "000011000011000000000",
    "000011000011010100000",
    "000011000011101000000",
    "000011000011111100000",
    "000011000100010000000",
    "000011000100100100000",
    "000011000100111000000",
    "000011000101001100000",
    "000011000101100000000",
    "000011000101110100000",
    "000011000110001000000",
    "000011000110011100000",
    "000011000110110000000",
    "000011000111000100000",
    "000011000111011000000",
    "000011000111101100000",
    "000011001000000000000",
    "000011001000010100000",
    "000011001000101000000",
    "000011001000111100000",
    "000011001001010000000",
    "000011001001100100000",
    "000011001001111000000",
    "000011001010001100000",
    "000011001010100000000",
    "000011001010110100000",
    "000011001011001000000",
    "000011001011011100000",
    "000011001011110000000",
    "000011001100000100000",
    "000011001100011000000",
    "000011001100101100000",
    "000011001101000000000",
    "000011001101010100000",
    "000011001101101000000",
    "000011001101111100000",
    "000011001110010000000",
    "000011001110100100000",
    "000011001110111000000",
    "000011001111001100000",
    "000011001111100000000",
    "000011001111110100000",
    "000011010000001000000",
    "000011010000011100000",
    "000011010000110000000",
    "000011010001000100000",
    "000011010001011000000",
    "000011010001101100000",
    "000011010010000000000",
    "000011010010010100000",
    "000011010010101000000",
    "000011010010111100000",
    "000011010011010000000",
    "000011010011100100000",
    "000011010011111000000",
    "000011010100001100000",
    "000011010100100000000",
    "000011010100110100000",
    "000011010101001000000",
    "000011010101011100000",
    "000011010101110000000",
    "000011010110000100000",
    "000011010110011000000",
    "000011010110101100000",
    "000011010111000000000",
    "000011010111010100000",
    "000011010111101000000",
    "000011010111111100000",
    "000011011000010000000",
    "000011011000100100000",
    "000011011000111000000",
    "000011011001001100000",
    "000011011001100000000",
    "000011011001110100000",
    "000011011010001000000",
    "000011011010011100000",
    "000011011010110000000",
    "000011011011000100000",
    "000011011011011000000",
    "000011011011101100000",
    "000011011100000000000",
    "000011011100010100000",
    "000011011100101000000",
    "000011011100111100000",
    "000011011101101110000",
    "000011100001000000000"
    );
    signal index : integer range 0 to 65535:= 0;
    signal count : std_logic_vector(20 downto 0):= (others => '0');
begin
    process(tempo_clock) begin
        if rising_edge(tempo_clock) then
            if reset_time = '0' then
                count <= count + 1;
                if count = time_ROM(index + 1) then
                    index <= index + 1;
                    checker_s <= '1';
                else 
                    checker_s <= '0';
                end if;     
            else
                index <= 0;
                checker_s <= '0';
                count <= (others => '0');
            end if;
        end if;
    end process;
    ROMaddress <= index;
end Behavioral;